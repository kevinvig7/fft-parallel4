`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.07.2019 14:35:16
// Design Name: 
// Module Name: BF
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module BF(
    input BFIn_up,
    input BFIn_down,
    output BFOut_up,
    output BFOut_down
    );
    
   
    
   assign  BFOut_up = BFIn_up;
    assign  BFOut_down = BFIn_down;
    
    
    
    
    
endmodule
